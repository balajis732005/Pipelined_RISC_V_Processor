module executeToMemory(
    input logic clock,
    input logic reset,
    input logic [31:0] pcAdderOut,
    input logic [31:0] aluOut,
    input logic isAluOutZero,
    
);



endmodule