module processor_tb;

    

endmodule