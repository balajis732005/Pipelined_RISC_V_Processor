module processor();
    
endmodule